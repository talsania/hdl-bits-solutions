module top_module (
    input [4:0] a, b, c, d, e, f,
    output [7:0] w, x, y, z );//
    wire [31:0] k;
    // assign { ... } = { ... };
    assign k={a,b,c,d,e,f,2'b11};
    assign w=k[31:24];
    assign x=k[23:16];
    assign y=k[15:8];
    assign z=k[7:0];
endmodule
