module top_module (
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);//
    wire x;
    wire [15:0] sum_lo, sum_hi;
    add16 instance1 (.a(a[15:0]),.b(b[15:0]),.cin(1'b0),.cout(x),.sum(sum_lo));
    add16 instance2 (.a(a[31:16]),.b(b[31:16]),.cin(x),.cout(),.sum(sum_hi));
    assign sum={sum_hi,sum_lo};
endmodule

module add1 ( input a, input b, input cin,   output sum, output cout );

// Full adder module here
    assign sum=a^b^cin;
    assign cout=a&b|a&cin|b&cin;
endmodule
